class cfg;
	static virtual intf vintf;
	static mailbox gen2drv=new();	
	static mailbox mon2cov=new();
	static mailbox mon2che=new();
endclass
