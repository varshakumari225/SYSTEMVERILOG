`include "mem.sv"
`include "c_intf.sv"
`include "mem_cfg.sv"
`include "mem_tx.sv"
`include "mem_gen.sv"
`include "mem_bfm.sv"
`include "monitor.sv"
`include "coverage.sv"
`include "checker.sv"
`include "mem_env.sv"
`include "test.sv"
`include "mem_top.sv"
